//-------------------------------------------------------------------------------------------------
module audio
//-------------------------------------------------------------------------------------------------
(
	input  wire      clock,
	input  wire      reset,
	input  wire[7:0] a,
	input  wire[7:0] b,
	input  wire[7:0] c,
	output wire[1:0] audio
);
//-------------------------------------------------------------------------------------------------

wire[9:0] ldacD = { 2'b00, a } + { 2'b00, b };
wire[9:0] rdacD = { 2'b00, b } + { 2'b00, c };

//-------------------------------------------------------------------------------------------------

dac #(.MSBI(9)) LDac
(
	.clock  (clock   ),
	.reset  (reset   ),
	.d      (ldacD   ),
	.q      (audio[0])
);

dac #(.MSBI(9)) RDac
(
	.clock  (clock   ),
	.reset  (reset   ),
	.d      (rdacD   ),
	.q      (audio[1])
);

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
